// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module cluster_clock_mux2
(
    input  logic clk0_i,
    input  logic clk1_i,
    input  logic clk_sel_i,
    output logic clk_o
  );

//  always_comb
//  begin
//    if (clk_sel_i == 1'b0)
//      clk_o = clk0_i;
//    else
//      clk_o = clk1_i;
//  end
   CKMUX2D0BWP12T clk_mux2 (
    .S(clk_sel_i),
    .I0(clk0_i),
    .I1(clk1_i),
    .Z(clk_o)
   );

endmodule
